module sys (
		input  wire  clk_clk,     //   clk.clk
		input  wire  reset_reset  // reset.reset
	);
endmodule

