// sys.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module sys (
		inout  wire [7:0] io_dq,               //              io.dq
		inout  wire       io_rwds,             //                .rwds
		output wire       io_ckout,            //                .ckout
		output wire       io_ckoutn,           //                .ckoutn
		output wire       io_csn,              //                .csn
		output wire       io_rstn,             //                .rstn
		output wire       jtag_uart_0_irq_irq, // jtag_uart_0_irq.irq
		input  wire       memrst_reset,        //          memrst.reset
		input  wire       refclk_clk,          //          refclk.clk
		input  wire       rst_reset            //             rst.reset
	);

	wire         hyperram_controller_0_coreclk_clk;                              // hyperram_controller_0:coreclk -> [intel_niosv_m_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:hyperram_controller_0_coreclk_clk, onchip_memory2_0:clk, rst_controller:clk, rst_controller_001:clk]
	wire  [31:0] intel_niosv_m_0_data_manager_readdata;                          // mm_interconnect_0:intel_niosv_m_0_data_manager_readdata -> intel_niosv_m_0:data_manager_readdata
	wire         intel_niosv_m_0_data_manager_waitrequest;                       // mm_interconnect_0:intel_niosv_m_0_data_manager_waitrequest -> intel_niosv_m_0:data_manager_waitrequest
	wire  [31:0] intel_niosv_m_0_data_manager_address;                           // intel_niosv_m_0:data_manager_address -> mm_interconnect_0:intel_niosv_m_0_data_manager_address
	wire         intel_niosv_m_0_data_manager_read;                              // intel_niosv_m_0:data_manager_read -> mm_interconnect_0:intel_niosv_m_0_data_manager_read
	wire   [3:0] intel_niosv_m_0_data_manager_byteenable;                        // intel_niosv_m_0:data_manager_byteenable -> mm_interconnect_0:intel_niosv_m_0_data_manager_byteenable
	wire         intel_niosv_m_0_data_manager_readdatavalid;                     // mm_interconnect_0:intel_niosv_m_0_data_manager_readdatavalid -> intel_niosv_m_0:data_manager_readdatavalid
	wire   [1:0] intel_niosv_m_0_data_manager_response;                          // mm_interconnect_0:intel_niosv_m_0_data_manager_response -> intel_niosv_m_0:data_manager_response
	wire         intel_niosv_m_0_data_manager_write;                             // intel_niosv_m_0:data_manager_write -> mm_interconnect_0:intel_niosv_m_0_data_manager_write
	wire  [31:0] intel_niosv_m_0_data_manager_writedata;                         // intel_niosv_m_0:data_manager_writedata -> mm_interconnect_0:intel_niosv_m_0_data_manager_writedata
	wire         intel_niosv_m_0_data_manager_writeresponsevalid;                // mm_interconnect_0:intel_niosv_m_0_data_manager_writeresponsevalid -> intel_niosv_m_0:data_manager_writeresponsevalid
	wire  [31:0] intel_niosv_m_0_instruction_manager_readdata;                   // mm_interconnect_0:intel_niosv_m_0_instruction_manager_readdata -> intel_niosv_m_0:instruction_manager_readdata
	wire         intel_niosv_m_0_instruction_manager_waitrequest;                // mm_interconnect_0:intel_niosv_m_0_instruction_manager_waitrequest -> intel_niosv_m_0:instruction_manager_waitrequest
	wire  [31:0] intel_niosv_m_0_instruction_manager_address;                    // intel_niosv_m_0:instruction_manager_address -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_address
	wire         intel_niosv_m_0_instruction_manager_read;                       // intel_niosv_m_0:instruction_manager_read -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_read
	wire         intel_niosv_m_0_instruction_manager_readdatavalid;              // mm_interconnect_0:intel_niosv_m_0_instruction_manager_readdatavalid -> intel_niosv_m_0:instruction_manager_readdatavalid
	wire   [1:0] intel_niosv_m_0_instruction_manager_response;                   // mm_interconnect_0:intel_niosv_m_0_instruction_manager_response -> intel_niosv_m_0:instruction_manager_response
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_csr_readdata;           // hyperram_controller_0:csr_readdata -> mm_interconnect_0:hyperram_controller_0_csr_readdata
	wire   [9:0] mm_interconnect_0_hyperram_controller_0_csr_address;            // mm_interconnect_0:hyperram_controller_0_csr_address -> hyperram_controller_0:csr_address
	wire         mm_interconnect_0_hyperram_controller_0_csr_read;               // mm_interconnect_0:hyperram_controller_0_csr_read -> hyperram_controller_0:csr_read
	wire         mm_interconnect_0_hyperram_controller_0_csr_readdatavalid;      // hyperram_controller_0:csr_readdatavalid -> mm_interconnect_0:hyperram_controller_0_csr_readdatavalid
	wire         mm_interconnect_0_hyperram_controller_0_csr_write;              // mm_interconnect_0:hyperram_controller_0_csr_write -> hyperram_controller_0:csr_write
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_csr_writedata;          // mm_interconnect_0:hyperram_controller_0_csr_writedata -> hyperram_controller_0:csr_writedata
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata;            // intel_niosv_m_0:dm_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest;         // intel_niosv_m_0:dm_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_address;             // mm_interconnect_0:intel_niosv_m_0_dm_agent_address -> intel_niosv_m_0:dm_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_read;                // mm_interconnect_0:intel_niosv_m_0_dm_agent_read -> intel_niosv_m_0:dm_agent_read
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid;       // intel_niosv_m_0:dm_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_write;               // mm_interconnect_0:intel_niosv_m_0_dm_agent_write -> intel_niosv_m_0:dm_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata;           // mm_interconnect_0:intel_niosv_m_0_dm_agent_writedata -> intel_niosv_m_0:dm_agent_writedata
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_s0_readdata;            // hyperram_controller_0:s0_readdata -> mm_interconnect_0:hyperram_controller_0_s0_readdata
	wire  [21:0] mm_interconnect_0_hyperram_controller_0_s0_address;             // mm_interconnect_0:hyperram_controller_0_s0_address -> hyperram_controller_0:s0_address
	wire         mm_interconnect_0_hyperram_controller_0_s0_read;                // mm_interconnect_0:hyperram_controller_0_s0_read -> hyperram_controller_0:s0_read
	wire         mm_interconnect_0_hyperram_controller_0_s0_readdatavalid;       // hyperram_controller_0:s0_readdatavalid -> mm_interconnect_0:hyperram_controller_0_s0_readdatavalid
	wire         mm_interconnect_0_hyperram_controller_0_s0_write;               // mm_interconnect_0:hyperram_controller_0_s0_write -> hyperram_controller_0:s0_write
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_s0_writedata;           // mm_interconnect_0:hyperram_controller_0_s0_writedata -> hyperram_controller_0:s0_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;               // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                 // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                  // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;               // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                    // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                    // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata;      // intel_niosv_m_0:timer_sw_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest;   // intel_niosv_m_0:timer_sw_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address;       // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_address -> intel_niosv_m_0:timer_sw_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read;          // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_read -> intel_niosv_m_0:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable;    // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_byteenable -> intel_niosv_m_0:timer_sw_agent_byteenable
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid; // intel_niosv_m_0:timer_sw_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write;         // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_write -> intel_niosv_m_0:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata;     // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_writedata -> intel_niosv_m_0:timer_sw_agent_writedata
	wire  [15:0] intel_niosv_m_0_platform_irq_rx_irq;                            // irq_mapper:sender_irq -> intel_niosv_m_0:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [intel_niosv_m_0:reset_reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:intel_niosv_m_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         hyperram_controller_0_corerst_reset;                            // hyperram_controller_0:corerst -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [mm_interconnect_0:hyperram_controller_0_csr_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:hyperram_controller_0_reset_controller_reset_bridge_in_reset_reset]

	hyperram_controller_top hyperram_controller_0 (
		.csr_address       (mm_interconnect_0_hyperram_controller_0_csr_address),       //              csr.address
		.csr_read          (mm_interconnect_0_hyperram_controller_0_csr_read),          //                 .read
		.csr_write         (mm_interconnect_0_hyperram_controller_0_csr_write),         //                 .write
		.csr_readdata      (mm_interconnect_0_hyperram_controller_0_csr_readdata),      //                 .readdata
		.csr_readdatavalid (mm_interconnect_0_hyperram_controller_0_csr_readdatavalid), //                 .readdatavalid
		.csr_writedata     (mm_interconnect_0_hyperram_controller_0_csr_writedata),     //                 .writedata
		.s0_address        (mm_interconnect_0_hyperram_controller_0_s0_address),        //               s0.address
		.s0_read           (mm_interconnect_0_hyperram_controller_0_s0_read),           //                 .read
		.s0_write          (mm_interconnect_0_hyperram_controller_0_s0_write),          //                 .write
		.s0_readdata       (mm_interconnect_0_hyperram_controller_0_s0_readdata),       //                 .readdata
		.s0_readdatavalid  (mm_interconnect_0_hyperram_controller_0_s0_readdatavalid),  //                 .readdatavalid
		.s0_writedata      (mm_interconnect_0_hyperram_controller_0_s0_writedata),      //                 .writedata
		.refclk            (refclk_clk),                                                //           refclk.clk
		.coreclk           (hyperram_controller_0_coreclk_clk),                         //          coreclk.clk
		.rst               (rst_reset),                                                 // reset_controller.reset
		.dq                (io_dq),                                                     //      hyperram_io.dq
		.rwds              (io_rwds),                                                   //                 .rwds
		.ckout             (io_ckout),                                                  //                 .ckout
		.ckoutn            (io_ckoutn),                                                 //                 .ckoutn
		.csn               (io_csn),                                                    //                 .csn
		.rstn              (io_rstn),                                                   //                 .rstn
		.memrst            (memrst_reset),                                              //     reset_memrst.reset
		.corerst           (hyperram_controller_0_corerst_reset)                        //          corerst.reset
	);

	sys_intel_niosv_m_0 intel_niosv_m_0 (
		.clk                               (hyperram_controller_0_coreclk_clk),                              //                 clk.clk
		.reset_reset                       (rst_controller_reset_out_reset),                                 //               reset.reset
		.platform_irq_rx_irq               (intel_niosv_m_0_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.timer_sw_agent_address            (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //      timer_sw_agent.address
		.timer_sw_agent_byteenable         (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_read               (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata           (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_write              (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //                    .write
		.timer_sw_agent_writedata          (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_waitrequest        (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //                    .waitrequest
		.timer_sw_agent_readdatavalid      (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.instruction_manager_readdata      (intel_niosv_m_0_instruction_manager_readdata),                   // instruction_manager.readdata
		.instruction_manager_waitrequest   (intel_niosv_m_0_instruction_manager_waitrequest),                //                    .waitrequest
		.instruction_manager_readdatavalid (intel_niosv_m_0_instruction_manager_readdatavalid),              //                    .readdatavalid
		.instruction_manager_response      (intel_niosv_m_0_instruction_manager_response),                   //                    .response
		.instruction_manager_address       (intel_niosv_m_0_instruction_manager_address),                    //                    .address
		.instruction_manager_read          (intel_niosv_m_0_instruction_manager_read),                       //                    .read
		.data_manager_readdata             (intel_niosv_m_0_data_manager_readdata),                          //        data_manager.readdata
		.data_manager_waitrequest          (intel_niosv_m_0_data_manager_waitrequest),                       //                    .waitrequest
		.data_manager_readdatavalid        (intel_niosv_m_0_data_manager_readdatavalid),                     //                    .readdatavalid
		.data_manager_response             (intel_niosv_m_0_data_manager_response),                          //                    .response
		.data_manager_address              (intel_niosv_m_0_data_manager_address),                           //                    .address
		.data_manager_read                 (intel_niosv_m_0_data_manager_read),                              //                    .read
		.data_manager_write                (intel_niosv_m_0_data_manager_write),                             //                    .write
		.data_manager_writedata            (intel_niosv_m_0_data_manager_writedata),                         //                    .writedata
		.data_manager_byteenable           (intel_niosv_m_0_data_manager_byteenable),                        //                    .byteenable
		.data_manager_writeresponsevalid   (intel_niosv_m_0_data_manager_writeresponsevalid),                //                    .writeresponsevalid
		.dm_agent_address                  (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //            dm_agent.address
		.dm_agent_read                     (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //                    .read
		.dm_agent_readdata                 (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //                    .readdata
		.dm_agent_write                    (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //                    .write
		.dm_agent_writedata                (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //                    .writedata
		.dm_agent_waitrequest              (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest),         //                    .waitrequest
		.dm_agent_readdatavalid            (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid)        //                    .readdatavalid
	);

	altera_avalon_jtag_uart #(
		.readBufferDepth            (64),
		.readIRQThreshold           (0),
		.useRegistersForReadBuffer  (0),
		.useRegistersForWriteBuffer (0),
		.writeBufferDepth           (64),
		.writeIRQThreshold          (0),
		.printingMethod             (0),
		.FIFO_WIDTH                 (8),
		.WR_WIDTHU                  (6),
		.RD_WIDTHU                  (6),
		.write_le                   ("ON"),
		.read_le                    ("ON"),
		.HEX_WRITE_DEPTH_STR        (64),
		.HEX_READ_DEPTH_STR         (64),
		.legacySignalAllow          (0)
	) jtag_uart_0 (
		.clk            (hyperram_controller_0_coreclk_clk),                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (jtag_uart_0_irq_irq)                                          //               irq.irq
	);

	sys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (hyperram_controller_0_coreclk_clk),                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	sys_mm_interconnect_0 mm_interconnect_0 (
		.hyperram_controller_0_coreclk_clk                                      (hyperram_controller_0_coreclk_clk),                              //                                    hyperram_controller_0_coreclk.clk
		.hyperram_controller_0_csr_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                             // hyperram_controller_0_csr_translator_reset_reset_bridge_in_reset.reset
		.hyperram_controller_0_reset_controller_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                             //     hyperram_controller_0_reset_controller_reset_bridge_in_reset.reset
		.intel_niosv_m_0_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),                                 //                      intel_niosv_m_0_reset_reset_bridge_in_reset.reset
		.intel_niosv_m_0_data_manager_address                                   (intel_niosv_m_0_data_manager_address),                           //                                     intel_niosv_m_0_data_manager.address
		.intel_niosv_m_0_data_manager_waitrequest                               (intel_niosv_m_0_data_manager_waitrequest),                       //                                                                 .waitrequest
		.intel_niosv_m_0_data_manager_byteenable                                (intel_niosv_m_0_data_manager_byteenable),                        //                                                                 .byteenable
		.intel_niosv_m_0_data_manager_read                                      (intel_niosv_m_0_data_manager_read),                              //                                                                 .read
		.intel_niosv_m_0_data_manager_readdata                                  (intel_niosv_m_0_data_manager_readdata),                          //                                                                 .readdata
		.intel_niosv_m_0_data_manager_readdatavalid                             (intel_niosv_m_0_data_manager_readdatavalid),                     //                                                                 .readdatavalid
		.intel_niosv_m_0_data_manager_write                                     (intel_niosv_m_0_data_manager_write),                             //                                                                 .write
		.intel_niosv_m_0_data_manager_writedata                                 (intel_niosv_m_0_data_manager_writedata),                         //                                                                 .writedata
		.intel_niosv_m_0_data_manager_response                                  (intel_niosv_m_0_data_manager_response),                          //                                                                 .response
		.intel_niosv_m_0_data_manager_writeresponsevalid                        (intel_niosv_m_0_data_manager_writeresponsevalid),                //                                                                 .writeresponsevalid
		.intel_niosv_m_0_instruction_manager_address                            (intel_niosv_m_0_instruction_manager_address),                    //                              intel_niosv_m_0_instruction_manager.address
		.intel_niosv_m_0_instruction_manager_waitrequest                        (intel_niosv_m_0_instruction_manager_waitrequest),                //                                                                 .waitrequest
		.intel_niosv_m_0_instruction_manager_read                               (intel_niosv_m_0_instruction_manager_read),                       //                                                                 .read
		.intel_niosv_m_0_instruction_manager_readdata                           (intel_niosv_m_0_instruction_manager_readdata),                   //                                                                 .readdata
		.intel_niosv_m_0_instruction_manager_readdatavalid                      (intel_niosv_m_0_instruction_manager_readdatavalid),              //                                                                 .readdatavalid
		.intel_niosv_m_0_instruction_manager_response                           (intel_niosv_m_0_instruction_manager_response),                   //                                                                 .response
		.hyperram_controller_0_csr_address                                      (mm_interconnect_0_hyperram_controller_0_csr_address),            //                                        hyperram_controller_0_csr.address
		.hyperram_controller_0_csr_write                                        (mm_interconnect_0_hyperram_controller_0_csr_write),              //                                                                 .write
		.hyperram_controller_0_csr_read                                         (mm_interconnect_0_hyperram_controller_0_csr_read),               //                                                                 .read
		.hyperram_controller_0_csr_readdata                                     (mm_interconnect_0_hyperram_controller_0_csr_readdata),           //                                                                 .readdata
		.hyperram_controller_0_csr_writedata                                    (mm_interconnect_0_hyperram_controller_0_csr_writedata),          //                                                                 .writedata
		.hyperram_controller_0_csr_readdatavalid                                (mm_interconnect_0_hyperram_controller_0_csr_readdatavalid),      //                                                                 .readdatavalid
		.hyperram_controller_0_s0_address                                       (mm_interconnect_0_hyperram_controller_0_s0_address),             //                                         hyperram_controller_0_s0.address
		.hyperram_controller_0_s0_write                                         (mm_interconnect_0_hyperram_controller_0_s0_write),               //                                                                 .write
		.hyperram_controller_0_s0_read                                          (mm_interconnect_0_hyperram_controller_0_s0_read),                //                                                                 .read
		.hyperram_controller_0_s0_readdata                                      (mm_interconnect_0_hyperram_controller_0_s0_readdata),            //                                                                 .readdata
		.hyperram_controller_0_s0_writedata                                     (mm_interconnect_0_hyperram_controller_0_s0_writedata),           //                                                                 .writedata
		.hyperram_controller_0_s0_readdatavalid                                 (mm_interconnect_0_hyperram_controller_0_s0_readdatavalid),       //                                                                 .readdatavalid
		.intel_niosv_m_0_dm_agent_address                                       (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //                                         intel_niosv_m_0_dm_agent.address
		.intel_niosv_m_0_dm_agent_write                                         (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //                                                                 .write
		.intel_niosv_m_0_dm_agent_read                                          (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //                                                                 .read
		.intel_niosv_m_0_dm_agent_readdata                                      (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //                                                                 .readdata
		.intel_niosv_m_0_dm_agent_writedata                                     (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //                                                                 .writedata
		.intel_niosv_m_0_dm_agent_readdatavalid                                 (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid),       //                                                                 .readdatavalid
		.intel_niosv_m_0_dm_agent_waitrequest                                   (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest),         //                                                                 .waitrequest
		.intel_niosv_m_0_timer_sw_agent_address                                 (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //                                   intel_niosv_m_0_timer_sw_agent.address
		.intel_niosv_m_0_timer_sw_agent_write                                   (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //                                                                 .write
		.intel_niosv_m_0_timer_sw_agent_read                                    (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //                                                                 .read
		.intel_niosv_m_0_timer_sw_agent_readdata                                (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //                                                                 .readdata
		.intel_niosv_m_0_timer_sw_agent_writedata                               (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //                                                                 .writedata
		.intel_niosv_m_0_timer_sw_agent_byteenable                              (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //                                                                 .byteenable
		.intel_niosv_m_0_timer_sw_agent_readdatavalid                           (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //                                                                 .readdatavalid
		.intel_niosv_m_0_timer_sw_agent_waitrequest                             (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //                                                                 .waitrequest
		.jtag_uart_0_avalon_jtag_slave_address                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),        //                                    jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),          //                                                                 .write
		.jtag_uart_0_avalon_jtag_slave_read                                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),           //                                                                 .read
		.jtag_uart_0_avalon_jtag_slave_readdata                                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),       //                                                                 .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),      //                                                                 .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),    //                                                                 .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),     //                                                                 .chipselect
		.onchip_memory2_0_s1_address                                            (mm_interconnect_0_onchip_memory2_0_s1_address),                  //                                              onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                              (mm_interconnect_0_onchip_memory2_0_s1_write),                    //                                                                 .write
		.onchip_memory2_0_s1_readdata                                           (mm_interconnect_0_onchip_memory2_0_s1_readdata),                 //                                                                 .readdata
		.onchip_memory2_0_s1_writedata                                          (mm_interconnect_0_onchip_memory2_0_s1_writedata),                //                                                                 .writedata
		.onchip_memory2_0_s1_byteenable                                         (mm_interconnect_0_onchip_memory2_0_s1_byteenable),               //                                                                 .byteenable
		.onchip_memory2_0_s1_chipselect                                         (mm_interconnect_0_onchip_memory2_0_s1_chipselect),               //                                                                 .chipselect
		.onchip_memory2_0_s1_clken                                              (mm_interconnect_0_onchip_memory2_0_s1_clken)                     //                                                                 .clken
	);

	sys_irq_mapper irq_mapper (
		.clk        (hyperram_controller_0_coreclk_clk),   //       clk.clk
		.reset      (rst_controller_reset_out_reset),      // clk_reset.reset
		.sender_irq (intel_niosv_m_0_platform_irq_rx_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (hyperram_controller_0_corerst_reset), // reset_in0.reset
		.clk            (hyperram_controller_0_coreclk_clk),   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (rst_reset),                          // reset_in0.reset
		.clk            (hyperram_controller_0_coreclk_clk),  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
