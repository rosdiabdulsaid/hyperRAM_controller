// sys_jamb.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module sys_jamb (
		input  wire       clk_clk,            //          clk.clk
		inout  wire [7:0] io_dq,              //           io.dq
		inout  wire       io_rwds,            //             .rwds
		output wire       io_ckout,           //             .ckout
		output wire       io_ckoutn,          //             .ckoutn
		output wire       io_csn,             //             .csn
		output wire       io_rstn,            //             .rstn
		output wire       master_reset_reset, // master_reset.reset
		input  wire       memrst_reset,       //       memrst.reset
		input  wire       reset_reset_n       //        reset.reset_n
	);

	wire         hyperram_controller_0_coreclk_clk;                         // hyperram_controller_0:coreclk -> [master_0:clk_clk, mm_interconnect_0:hyperram_controller_0_coreclk_clk, rst_controller:clk, rst_controller_001:clk]
	wire         hyperram_controller_0_corerst_reset;                       // hyperram_controller_0:corerst -> [master_0:clk_reset_reset, rst_controller_001:reset_in0]
	wire  [31:0] master_0_master_readdata;                                  // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                               // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                   // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                      // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                             // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                     // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                 // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_csr_readdata;      // hyperram_controller_0:csr_readdata -> mm_interconnect_0:hyperram_controller_0_csr_readdata
	wire         mm_interconnect_0_hyperram_controller_0_csr_waitrequest;   // hyperram_controller_0:csr_waitrequest -> mm_interconnect_0:hyperram_controller_0_csr_waitrequest
	wire   [9:0] mm_interconnect_0_hyperram_controller_0_csr_address;       // mm_interconnect_0:hyperram_controller_0_csr_address -> hyperram_controller_0:csr_address
	wire         mm_interconnect_0_hyperram_controller_0_csr_read;          // mm_interconnect_0:hyperram_controller_0_csr_read -> hyperram_controller_0:csr_read
	wire         mm_interconnect_0_hyperram_controller_0_csr_readdatavalid; // hyperram_controller_0:csr_readdatavalid -> mm_interconnect_0:hyperram_controller_0_csr_readdatavalid
	wire         mm_interconnect_0_hyperram_controller_0_csr_write;         // mm_interconnect_0:hyperram_controller_0_csr_write -> hyperram_controller_0:csr_write
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_csr_writedata;     // mm_interconnect_0:hyperram_controller_0_csr_writedata -> hyperram_controller_0:csr_writedata
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_s0_readdata;       // hyperram_controller_0:s0_readdata -> mm_interconnect_0:hyperram_controller_0_s0_readdata
	wire         mm_interconnect_0_hyperram_controller_0_s0_waitrequest;    // hyperram_controller_0:s0_waitrequest -> mm_interconnect_0:hyperram_controller_0_s0_waitrequest
	wire  [21:0] mm_interconnect_0_hyperram_controller_0_s0_address;        // mm_interconnect_0:hyperram_controller_0_s0_address -> hyperram_controller_0:s0_address
	wire         mm_interconnect_0_hyperram_controller_0_s0_read;           // mm_interconnect_0:hyperram_controller_0_s0_read -> hyperram_controller_0:s0_read
	wire         mm_interconnect_0_hyperram_controller_0_s0_readdatavalid;  // hyperram_controller_0:s0_readdatavalid -> mm_interconnect_0:hyperram_controller_0_s0_readdatavalid
	wire         mm_interconnect_0_hyperram_controller_0_s0_write;          // mm_interconnect_0:hyperram_controller_0_s0_write -> hyperram_controller_0:s0_write
	wire  [31:0] mm_interconnect_0_hyperram_controller_0_s0_writedata;      // mm_interconnect_0:hyperram_controller_0_s0_writedata -> hyperram_controller_0:s0_writedata
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [mm_interconnect_0:hyperram_controller_0_csr_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:hyperram_controller_0_reset_controller_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_master_translator_reset_reset_bridge_in_reset_reset]

	hyperram_controller_top hyperram_controller_0 (
		.csr_address       (mm_interconnect_0_hyperram_controller_0_csr_address),       //              csr.address
		.csr_read          (mm_interconnect_0_hyperram_controller_0_csr_read),          //                 .read
		.csr_write         (mm_interconnect_0_hyperram_controller_0_csr_write),         //                 .write
		.csr_readdata      (mm_interconnect_0_hyperram_controller_0_csr_readdata),      //                 .readdata
		.csr_readdatavalid (mm_interconnect_0_hyperram_controller_0_csr_readdatavalid), //                 .readdatavalid
		.csr_writedata     (mm_interconnect_0_hyperram_controller_0_csr_writedata),     //                 .writedata
		.csr_waitrequest   (mm_interconnect_0_hyperram_controller_0_csr_waitrequest),   //                 .waitrequest
		.s0_address        (mm_interconnect_0_hyperram_controller_0_s0_address),        //               s0.address
		.s0_read           (mm_interconnect_0_hyperram_controller_0_s0_read),           //                 .read
		.s0_write          (mm_interconnect_0_hyperram_controller_0_s0_write),          //                 .write
		.s0_readdata       (mm_interconnect_0_hyperram_controller_0_s0_readdata),       //                 .readdata
		.s0_readdatavalid  (mm_interconnect_0_hyperram_controller_0_s0_readdatavalid),  //                 .readdatavalid
		.s0_writedata      (mm_interconnect_0_hyperram_controller_0_s0_writedata),      //                 .writedata
		.s0_waitrequest    (mm_interconnect_0_hyperram_controller_0_s0_waitrequest),    //                 .waitrequest
		.refclk            (clk_clk),                                                   //           refclk.clk
		.coreclk           (hyperram_controller_0_coreclk_clk),                         //          coreclk.clk
		.rst               (~reset_reset_n),                                            // reset_controller.reset
		.dq                (io_dq),                                                     //      hyperram_io.dq
		.rwds              (io_rwds),                                                   //                 .rwds
		.ckout             (io_ckout),                                                  //                 .ckout
		.ckoutn            (io_ckoutn),                                                 //                 .ckoutn
		.csn               (io_csn),                                                    //                 .csn
		.rstn              (io_rstn),                                                   //                 .rstn
		.corerst           (hyperram_controller_0_corerst_reset),                       //          corerst.reset
		.memrst            (memrst_reset)                                               //     reset_memrst.reset
	);

	sys_jamb_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (hyperram_controller_0_coreclk_clk),   //          clk.clk
		.clk_reset_reset      (hyperram_controller_0_corerst_reset), //    clk_reset.reset
		.master_address       (master_0_master_address),             //       master.address
		.master_readdata      (master_0_master_readdata),            //             .readdata
		.master_read          (master_0_master_read),                //             .read
		.master_write         (master_0_master_write),               //             .write
		.master_writedata     (master_0_master_writedata),           //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),         //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid),       //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),          //             .byteenable
		.master_reset_reset   (master_reset_reset)                   // master_reset.reset
	);

	sys_jamb_mm_interconnect_0 mm_interconnect_0 (
		.hyperram_controller_0_coreclk_clk                                      (hyperram_controller_0_coreclk_clk),                         //                                    hyperram_controller_0_coreclk.clk
		.hyperram_controller_0_csr_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // hyperram_controller_0_csr_translator_reset_reset_bridge_in_reset.reset
		.hyperram_controller_0_reset_controller_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                            //     hyperram_controller_0_reset_controller_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset                         (rst_controller_001_reset_out_reset),                        //                         master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_translator_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                        //           master_0_master_translator_reset_reset_bridge_in_reset.reset
		.master_0_master_address                                                (master_0_master_address),                                   //                                                  master_0_master.address
		.master_0_master_waitrequest                                            (master_0_master_waitrequest),                               //                                                                 .waitrequest
		.master_0_master_byteenable                                             (master_0_master_byteenable),                                //                                                                 .byteenable
		.master_0_master_read                                                   (master_0_master_read),                                      //                                                                 .read
		.master_0_master_readdata                                               (master_0_master_readdata),                                  //                                                                 .readdata
		.master_0_master_readdatavalid                                          (master_0_master_readdatavalid),                             //                                                                 .readdatavalid
		.master_0_master_write                                                  (master_0_master_write),                                     //                                                                 .write
		.master_0_master_writedata                                              (master_0_master_writedata),                                 //                                                                 .writedata
		.hyperram_controller_0_csr_address                                      (mm_interconnect_0_hyperram_controller_0_csr_address),       //                                        hyperram_controller_0_csr.address
		.hyperram_controller_0_csr_write                                        (mm_interconnect_0_hyperram_controller_0_csr_write),         //                                                                 .write
		.hyperram_controller_0_csr_read                                         (mm_interconnect_0_hyperram_controller_0_csr_read),          //                                                                 .read
		.hyperram_controller_0_csr_readdata                                     (mm_interconnect_0_hyperram_controller_0_csr_readdata),      //                                                                 .readdata
		.hyperram_controller_0_csr_writedata                                    (mm_interconnect_0_hyperram_controller_0_csr_writedata),     //                                                                 .writedata
		.hyperram_controller_0_csr_readdatavalid                                (mm_interconnect_0_hyperram_controller_0_csr_readdatavalid), //                                                                 .readdatavalid
		.hyperram_controller_0_csr_waitrequest                                  (mm_interconnect_0_hyperram_controller_0_csr_waitrequest),   //                                                                 .waitrequest
		.hyperram_controller_0_s0_address                                       (mm_interconnect_0_hyperram_controller_0_s0_address),        //                                         hyperram_controller_0_s0.address
		.hyperram_controller_0_s0_write                                         (mm_interconnect_0_hyperram_controller_0_s0_write),          //                                                                 .write
		.hyperram_controller_0_s0_read                                          (mm_interconnect_0_hyperram_controller_0_s0_read),           //                                                                 .read
		.hyperram_controller_0_s0_readdata                                      (mm_interconnect_0_hyperram_controller_0_s0_readdata),       //                                                                 .readdata
		.hyperram_controller_0_s0_writedata                                     (mm_interconnect_0_hyperram_controller_0_s0_writedata),      //                                                                 .writedata
		.hyperram_controller_0_s0_readdatavalid                                 (mm_interconnect_0_hyperram_controller_0_s0_readdatavalid),  //                                                                 .readdatavalid
		.hyperram_controller_0_s0_waitrequest                                   (mm_interconnect_0_hyperram_controller_0_s0_waitrequest)     //                                                                 .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.clk            (hyperram_controller_0_coreclk_clk), //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_in1      (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (hyperram_controller_0_corerst_reset), // reset_in0.reset
		.clk            (hyperram_controller_0_coreclk_clk),   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
